--- This is the working code of a Descriptor Bypass Controller for the XDMA IP from Xilinx. 
--References : https://github.com/rsarwar87/xdma_dsc_byp_cltr

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity desc_byp is
generic(

--User Parameters
 
S_AXI_DATA_WIDTH : integer := 32;
S_AXI_ADDR_WIDTH : integer := 5
);

--  Ports

port(
                dsc_byp_ctl         : out std_logic_vector (15 downto 0);
                dsc_byp_dst_addr    : out std_logic_vector (63 downto 0);
                dsc_byp_src_addr    : out std_logic_vector (63 downto 0);
                dsc_byp_length      : out std_logic_vector (27 downto 0);
                dsc_byp_ready       : in  std_logic;
                dsc_byp_load        : out std_logic;

-- User ports ends
-- Do not modify the ports beyond this line

-- Global Clock Signal
S_AXI_ACLK : in std_logic;
-- Global Reset Signal. This Signal is Active LOW
S_AXI_ARESETN : in std_logic;
-- Write address (issued by master, acceped by Slave)
S_AXI_AWADDR : in std_logic_vector(S_AXI_ADDR_WIDTH-1 downto 0);
-- Write channel Protection type. This signal indicates the
    -- privilege and security level of the transaction, and whether
    -- the transaction is a data access or an instruction access.
S_AXI_AWPROT : in std_logic_vector(2 downto 0);
-- Write address valid. This signal indicates that the master signaling
    -- valid write address and control information.
S_AXI_AWVALID : in std_logic;
-- Write address ready. This signal indicates that the slave is ready
    -- to accept an address and associated control signals.
S_AXI_AWREADY : out std_logic;
-- Write data (issued by master, acceped by Slave)
S_AXI_WDATA : in std_logic_vector(S_AXI_DATA_WIDTH-1 downto 0);
-- Write strobes. This signal indicates which byte lanes hold
    -- valid data. There is one write strobe bit for each eight
    -- bits of the write data bus.    
S_AXI_WSTRB : in std_logic_vector((S_AXI_DATA_WIDTH/8)-1 downto 0);
-- Write valid. This signal indicates that valid write
    -- data and strobes are available.
S_AXI_WVALID : in std_logic;
-- Write ready. This signal indicates that the slave
    -- can accept the write data.
S_AXI_WREADY : out std_logic;
-- Write response. This signal indicates the status
    -- of the write transaction.
S_AXI_BRESP : out std_logic_vector(1 downto 0);
-- Write response valid. This signal indicates that the channel
    -- is signaling a valid write response.
S_AXI_BVALID : out std_logic;
-- Response ready. This signal indicates that the master
    -- can accept a write response.
S_AXI_BREADY : in std_logic;
-- Read address (issued by master, acceped by Slave)
S_AXI_ARADDR : in std_logic_vector(S_AXI_ADDR_WIDTH-1 downto 0);
-- Protection type. This signal indicates the privilege
    -- and security level of the transaction, and whether the
    -- transaction is a data access or an instruction access.
S_AXI_ARPROT : in std_logic_vector(2 downto 0);
-- Read address valid. This signal indicates that the channel
    -- is signaling valid read address and control information.
S_AXI_ARVALID : in std_logic;
-- Read address ready. This signal indicates that the slave is
    -- ready to accept an address and associated control signals.
S_AXI_ARREADY : out std_logic;
-- Read data (issued by slave)
S_AXI_RDATA : out std_logic_vector(S_AXI_DATA_WIDTH-1 downto 0);
-- Read response. This signal indicates the status of the
    -- read transfer.
S_AXI_RRESP : out std_logic_vector(1 downto 0);
-- Read valid. This signal indicates that the channel is
    -- signaling the required read data.
S_AXI_RVALID : out std_logic;
-- Read ready. This signal indicates that the master can
    -- accept the read data and response information.
S_AXI_RREADY : in std_logic
);
end desc_byp;
architecture arch_imp of desc_byp is

-- AXI4LITE signals
signal axi_awaddr : std_logic_vector(S_AXI_ADDR_WIDTH-1 downto 0);
signal axi_awready : std_logic;
signal axi_wready : std_logic;
signal axi_bresp : std_logic_vector(1 downto 0);
signal axi_bvalid : std_logic;
signal axi_araddr : std_logic_vector(S_AXI_ADDR_WIDTH-1 downto 0);
signal axi_arready : std_logic;
signal axi_rdata : std_logic_vector(S_AXI_DATA_WIDTH-1 downto 0);
signal axi_rresp : std_logic_vector(1 downto 0);
signal axi_rvalid : std_logic;

-- Example-specific design signals
-- local parameter for addressing 32 bit / 64 bit S_AXI_DATA_WIDTH
-- ADDR_LSB is used for addressing 32/64 bit registers/memories
-- ADDR_LSB = 2 for 32 bits (n downto 2)
-- ADDR_LSB = 3 for 64 bits (n downto 3)
constant ADDR_LSB  : integer := (S_AXI_DATA_WIDTH/32)+ 1;
constant OPT_MEM_ADDR_BITS : integer := 2;
------------------------------------------------
---- Signals for user logic register space example
--------------------------------------------------
---- Number of Slave Registers 8
signal slv_reg0 :std_logic_vector(S_AXI_DATA_WIDTH-1 downto 0);
signal slv_reg1 :std_logic_vector(S_AXI_DATA_WIDTH-1 downto 0);
signal slv_reg2 :std_logic_vector(S_AXI_DATA_WIDTH-1 downto 0);
signal slv_reg3 :std_logic_vector(S_AXI_DATA_WIDTH-1 downto 0);
signal slv_reg4 :std_logic_vector(S_AXI_DATA_WIDTH-1 downto 0);
signal slv_reg5 :std_logic_vector(S_AXI_DATA_WIDTH-1 downto 0);
signal slv_reg6 :std_logic_vector(S_AXI_DATA_WIDTH-1 downto 0);
signal slv_reg7 :std_logic_vector(S_AXI_DATA_WIDTH-1 downto 0);
signal slv_reg_rden : std_logic;
signal slv_reg_wren : std_logic;
signal reg_data_out :std_logic_vector(S_AXI_DATA_WIDTH-1 downto 0);
signal byte_index : integer;
signal aw_en : std_logic;

    signal bypass_ctl          : std_logic_vector (15 downto 0) := (others => '0');
    signal bypass_dst_addr     : std_logic_vector (63 downto 0) := (others => '0');
    signal bypass_src_addr     : std_logic_vector (63 downto 0) := (others => '0');
    signal bypass_length       : std_logic_vector (27 downto 0) := (others => '0');
    signal bypass_start        : std_logic := '0';
    signal bypass_reset        : std_logic := '0';
    signal bypass_cyclic       : std_logic := '0';
    signal bypass_repeat       : std_logic_vector (31 downto 0) := (others => '0');
    signal bypass_count        : std_logic_vector (30 downto 0) := (others => '0');
    signal bypass_busy         : std_logic := '0';
    signal bypass_awk          : std_logic := '0';
    signal bypass_src_mm, bypass_dst_mm : std_logic := '0';
    signal bypass_addr_cnt     : std_logic_vector (63 downto 0) := (others => '0');
   
begin  
-- I/O Connections assignments
-- Control For the XDMA Control Interface
        bypass_ctl <= slv_reg0(15 downto 0);
-- Destination Address in the Card/Host for the DMA transfer
        bypass_dst_addr <= slv_reg1 & slv_reg2;
-- Source Address of the Host/Card for the DMA transfer
        bypass_src_addr <= slv_reg3 & slv_reg4;
-- Length of the DMA transfer
        bypass_length <= slv_reg5(27 downto 0);
-- Reset the whole controller
        bypass_reset <= slv_reg7(31);
-- Set if Destination is memory mapped. Clear if it is streaming
        bypass_dst_mm <= slv_reg7(3);
-- Set if Source is memory mapped. Clear if it is streaming
        bypass_src_mm <= slv_reg7(2);
-- Loop the Controller's operations
        bypass_cyclic <= slv_reg7(1);
-- Start feeding the values to the Descriptor Bypass ports
        bypass_start <= slv_reg7(0);
-- Repeat the controller's operations 'n' times. Where n is the number you give to the register
        bypass_repeat <= slv_reg6;

S_AXI_AWREADY <= axi_awready;
S_AXI_WREADY <= axi_wready;
S_AXI_BRESP <= axi_bresp;
S_AXI_BVALID <= axi_bvalid;
S_AXI_ARREADY <= axi_arready;
S_AXI_RDATA <= axi_rdata;
S_AXI_RRESP <= axi_rresp;
S_AXI_RVALID <= axi_rvalid;
-- Implement axi_awready generation
-- axi_awready is asserted for one S_AXI_ACLK clock cycle when both
-- S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_awready is
-- de-asserted when reset is low.

process (S_AXI_ACLK)
begin
 if rising_edge(S_AXI_ACLK) then
   if S_AXI_ARESETN = '0' then
     axi_awready <= '0';
     aw_en <= '1';
   else
     if (axi_awready = '0' and S_AXI_AWVALID = '1' and S_AXI_WVALID = '1' and aw_en = '1') then
       -- slave is ready to accept write address when
       -- there is a valid write address and write data
       -- on the write address and data bus. This design
       -- expects no outstanding transactions.
       axi_awready <= '1';
       elsif (S_AXI_BREADY = '1' and axi_bvalid = '1') then
           aw_en <= '1';
        axi_awready <= '0';
     else
       axi_awready <= '0';
     end if;
   end if;
 end if;
end process;

-- Implement axi_awaddr latching
-- This process is used to latch the address when both
-- S_AXI_AWVALID and S_AXI_WVALID are valid.

process (S_AXI_ACLK)
begin
 if rising_edge(S_AXI_ACLK) then
   if S_AXI_ARESETN = '0' then
     axi_awaddr <= (others => '0');
   else
     if (axi_awready = '0' and S_AXI_AWVALID = '1' and S_AXI_WVALID = '1' and aw_en = '1') then
       -- Write Address latching
       axi_awaddr <= S_AXI_AWADDR;
     end if;
   end if;
 end if;                  
end process;

-- Implement axi_wready generation
-- axi_wready is asserted for one S_AXI_ACLK clock cycle when both
-- S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_wready is
-- de-asserted when reset is low.

process (S_AXI_ACLK)
begin
 if rising_edge(S_AXI_ACLK) then
   if S_AXI_ARESETN = '0' then
     axi_wready <= '0';
   else
     if (axi_wready = '0' and S_AXI_WVALID = '1' and S_AXI_AWVALID = '1' and aw_en = '1') then
         -- slave is ready to accept write data when
         -- there is a valid write address and write data
         -- on the write address and data bus. This design
         -- expects no outstanding transactions.          
         axi_wready <= '1';
     else
       axi_wready <= '0';
     end if;
   end if;
 end if;
end process;

-- Implement memory mapped register select and write logic generation
-- The write data is accepted and written to memory mapped registers when
-- axi_awready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted. Write strobes are used to
-- select byte enables of slave registers while writing.
-- These registers are cleared when reset (active low) is applied.
-- Slave register write enable is asserted when valid address and data are available
-- and the slave is ready to accept the write address and write data.
slv_reg_wren <= axi_wready and S_AXI_WVALID and axi_awready and S_AXI_AWVALID ;

process (S_AXI_ACLK)
variable loc_addr :std_logic_vector(OPT_MEM_ADDR_BITS downto 0);
begin
 if rising_edge(S_AXI_ACLK) then
   if S_AXI_ARESETN = '0' then
     slv_reg0 <= (others => '0');
     slv_reg1 <= (others => '0');
     slv_reg2 <= (others => '0');
     slv_reg3 <= (others => '0');
     slv_reg4 <= (others => '0');
     slv_reg5 <= (others => '0');
     slv_reg6 <= (others => '0');
     slv_reg7 <= (others => '0');
   else
     loc_addr := axi_awaddr(ADDR_LSB + OPT_MEM_ADDR_BITS downto ADDR_LSB);
     if (slv_reg_wren = '1') then
       case loc_addr is
         when b"000" =>
           for byte_index in 0 to (S_AXI_DATA_WIDTH/8-1) loop
             if ( S_AXI_WSTRB(byte_index) = '1' ) then
               -- Respective byte enables are asserted as per write strobes                  
               -- slave registor 0
               slv_reg0(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
             end if;
           end loop;
         when b"001" =>
           for byte_index in 0 to (S_AXI_DATA_WIDTH/8-1) loop
             if ( S_AXI_WSTRB(byte_index) = '1' ) then
               -- Respective byte enables are asserted as per write strobes                  
               -- slave registor 1
               slv_reg1(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
             end if;
           end loop;
         when b"010" =>
           for byte_index in 0 to (S_AXI_DATA_WIDTH/8-1) loop
             if ( S_AXI_WSTRB(byte_index) = '1' ) then
               -- Respective byte enables are asserted as per write strobes                  
               -- slave registor 2
               slv_reg2(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
             end if;
           end loop;
         when b"011" =>
           for byte_index in 0 to (S_AXI_DATA_WIDTH/8-1) loop
             if ( S_AXI_WSTRB(byte_index) = '1' ) then
               -- Respective byte enables are asserted as per write strobes                  
               -- slave registor 3
               slv_reg3(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
             end if;
           end loop;
         when b"100" =>
           for byte_index in 0 to (S_AXI_DATA_WIDTH/8-1) loop
             if ( S_AXI_WSTRB(byte_index) = '1' ) then
               -- Respective byte enables are asserted as per write strobes                  
               -- slave registor 4
               slv_reg4(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
             end if;
           end loop;
         when b"101" =>
           for byte_index in 0 to (S_AXI_DATA_WIDTH/8-1) loop
             if ( S_AXI_WSTRB(byte_index) = '1' ) then
               -- Respective byte enables are asserted as per write strobes                  
               -- slave registor 5
               slv_reg5(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
             end if;
           end loop;
         when b"110" =>
           for byte_index in 0 to (S_AXI_DATA_WIDTH/8-1) loop
             if ( S_AXI_WSTRB(byte_index) = '1' ) then
               -- Respective byte enables are asserted as per write strobes                  
               -- slave registor 6
               slv_reg6(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
             end if;
           end loop;
         when b"111" =>
           for byte_index in 0 to (S_AXI_DATA_WIDTH/8-1) loop
             if ( S_AXI_WSTRB(byte_index) = '1' ) then
               -- Respective byte enables are asserted as per write strobes                  
               -- slave registor 7
               slv_reg7(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
             end if;
           end loop;
         when others =>
           slv_reg0 <= slv_reg0;
           slv_reg1 <= slv_reg1;
           slv_reg2 <= slv_reg2;
           slv_reg3 <= slv_reg3;
           slv_reg4 <= slv_reg4;
           slv_reg5 <= slv_reg5;
           slv_reg6 <= slv_reg6;
           slv_reg7 <= slv_reg7;
                   
       end case;
     end if;
     if (bypass_awk = '1') then
              slv_reg7(0) <= '0';
          end if;
   end if;
 end if;                  
end process;

-- Implement write response logic generation
-- The write response and response valid signals are asserted by the slave
-- when axi_wready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted.  
-- This marks the acceptance of address and indicates the status of
-- write transaction.

process (S_AXI_ACLK)
begin
 if rising_edge(S_AXI_ACLK) then
   if S_AXI_ARESETN = '0' then
     axi_bvalid  <= '0';
     axi_bresp   <= "00"; --need to work more on the responses
   else
     if (axi_awready = '1' and S_AXI_AWVALID = '1' and axi_wready = '1' and S_AXI_WVALID = '1' and axi_bvalid = '0'  ) then
       axi_bvalid <= '1';
       axi_bresp  <= "00";
     elsif (S_AXI_BREADY = '1' and axi_bvalid = '1') then   --check if bready is asserted while bvalid is high)
       axi_bvalid <= '0';                                 -- (there is a possibility that bready is always asserted high)
     end if;
   end if;
 end if;                  
end process;

-- Implement axi_arready generation
-- axi_arready is asserted for one S_AXI_ACLK clock cycle when
-- S_AXI_ARVALID is asserted. axi_awready is
-- de-asserted when reset (active low) is asserted.
-- The read address is also latched when S_AXI_ARVALID is
-- asserted. axi_araddr is reset to zero on reset assertion.

process (S_AXI_ACLK)
begin
 if rising_edge(S_AXI_ACLK) then
   if S_AXI_ARESETN = '0' then
     axi_arready <= '0';
     axi_araddr  <= (others => '1');
   else
     if (axi_arready = '0' and S_AXI_ARVALID = '1') then
       -- indicates that the slave has acceped the valid read address
       axi_arready <= '1';
       -- Read Address latching
       axi_araddr  <= S_AXI_ARADDR;          
     else
       axi_arready <= '0';
     end if;
   end if;
 end if;                  
end process;

-- Implement axi_arvalid generation
-- axi_rvalid is asserted for one S_AXI_ACLK clock cycle when both
-- S_AXI_ARVALID and axi_arready are asserted. The slave registers
-- data are available on the axi_rdata bus at this instance. The
-- assertion of axi_rvalid marks the validity of read data on the
-- bus and axi_rresp indicates the status of read transaction.axi_rvalid
-- is deasserted on reset (active low). axi_rresp and axi_rdata are
-- cleared to zero on reset (active low).  
process (S_AXI_ACLK)
begin
 if rising_edge(S_AXI_ACLK) then
   if S_AXI_ARESETN = '0' then
     axi_rvalid <= '0';
     axi_rresp  <= "00";
   else
     if (axi_arready = '1' and S_AXI_ARVALID = '1' and axi_rvalid = '0') then
       -- Valid read data is available at the read data bus
       axi_rvalid <= '1';
       axi_rresp  <= "00"; -- 'OKAY' response
     elsif (axi_rvalid = '1' and S_AXI_RREADY = '1') then
       -- Read data is accepted by the master
       axi_rvalid <= '0';
     end if;            
   end if;
 end if;
end process;

-- Implement memory mapped register select and read logic generation
-- Slave register read enable is asserted when valid address is available
-- and the slave is ready to accept the read address.

slv_reg_rden <= axi_arready and S_AXI_ARVALID and (not axi_rvalid) ;

process (slv_reg0, slv_reg1, slv_reg2, slv_reg3, slv_reg4, slv_reg5, slv_reg6, slv_reg7, axi_araddr, S_AXI_ARESETN, slv_reg_rden)
variable loc_addr :std_logic_vector(OPT_MEM_ADDR_BITS downto 0);
begin
   -- Address decoding for reading registers
   loc_addr := axi_araddr(ADDR_LSB + OPT_MEM_ADDR_BITS downto ADDR_LSB);
   case loc_addr is
     when b"000" =>
       reg_data_out <= slv_reg0;
     when b"001" =>
       reg_data_out <= slv_reg1;
     when b"010" =>
       reg_data_out <= slv_reg2;
     when b"011" =>
       reg_data_out <= slv_reg3;
     when b"100" =>
       reg_data_out <= slv_reg4;
     when b"101" =>
       reg_data_out <= slv_reg5;
     when b"110" =>
       reg_data_out <= slv_reg6;
     when b"111" =>
       reg_data_out <= slv_reg7;
     when others =>
       reg_data_out  <= (others => '0');
   end case;
end process;

-- Output register or memory read data

process( S_AXI_ACLK ) is
begin
 if (rising_edge (S_AXI_ACLK)) then
   if ( S_AXI_ARESETN = '0' ) then
     axi_rdata  <= (others => '0');
   else
     if (slv_reg_rden = '1') then
       -- When there is a valid read address (S_AXI_ARVALID) with
       -- acceptance of read address by the slave (axi_arready),
       -- output the read dada
       -- Read address mux
         axi_rdata <= reg_data_out;     -- register read data
     end if;  
   end if;
 end if;
end process;
   
    -- Output of the Descriptor Bypass Ports
   
    process(S_AXI_ACLK, S_AXI_ARESETN) is
   variable cnt : integer := 4;
    begin
        if (S_AXI_ARESETN = '0') then
            cnt := 1;
            dsc_byp_load <= '0';
            dsc_byp_ctl <= (others => '0');
            dsc_byp_src_addr <= (others => '0');
            dsc_byp_dst_addr <= (others => '0');
            dsc_byp_length <= (others => '0');
            bypass_count <= (others => '0');
            bypass_addr_cnt <= (others => '0');
        elsif (rising_edge(S_AXI_ACLK)) then
                if (dsc_byp_ready = '1') then
                    if (cnt = 0) then
                        cnt := 1;
                        dsc_byp_ctl <= bypass_ctl;
                        if (bypass_src_mm = '0') then
                            dsc_byp_src_addr <= bypass_src_addr;
                        else
                            dsc_byp_src_addr <= std_logic_vector(unsigned(bypass_src_addr));
                            --dsc_byp_src_addr <= std_logic_vector(unsigned(bypass_src_addr) + unsigned(bypass_addr_cnt));
                        end if;
                        if (bypass_dst_mm = '1') then
                            --dsc_byp_dst_addr <= std_logic_vector(unsigned(bypass_dst_addr) + unsigned(bypass_addr_cnt));
                            dsc_byp_dst_addr <= std_logic_vector(unsigned(bypass_dst_addr));
                        else
                            dsc_byp_dst_addr <= bypass_dst_addr;
                        end if;
                        dsc_byp_length <= bypass_length;
                        --bypass_addr_cnt <= std_logic_vector(unsigned(bypass_addr_cnt) + unsigned(bypass_length));
                        dsc_byp_load <= '1';
                        --bypass_count <= std_logic_vector(unsigned(bypass_count) + 1);
                        --byp_addr_cnt <= (others => '0');
                    else 
                        dsc_byp_load <= '0';
                        cnt := cnt - 1;
                        --if (bypass_repeat = bypass_count) then 
                            --bypass_count <= (others => '0');
                            --bypass_addr_cnt <= (others => '0');
                        --end if;
                    end if;
                else
                    cnt := 1;
                end if;
        end if;
    end process;
 
   
end arch_imp;

